module top(
    input clk,
    input reset,
    input cont,
    input run,
    output [7:0] an,
    output [6:0] seg,
    output dp,
    output [15:0] led
);

    

endmodule // top